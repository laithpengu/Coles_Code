/*
 *
 *   File Name:    cpu.sv
 *   Date Created: Mon May 01 2023
 *   Author:       Cole Cavanagh
 *   Description:  Control Logic for 316 HW 5
 *
 */

module cpu(


);

endmodule